module verilator_warning;
   reg val;
endmodule
