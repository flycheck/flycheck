module verilog_verilator_warning;
   reg val;
endmodule
