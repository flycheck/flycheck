entity syntax_error is
end entity syntax_error

